`ifndef CONST
`define CONST

// The instruction segments
`define FUNCT2  31:30
`define RS2     24:20    
`define SHAMT   24:20
`define RS1     19:15
`define FUNCT   14:12
`define RD      11:7
`define OP      6:0

// Define your own constants here, for use in the processor!

`endif //CONST
